// *********************************************************************************
// Project Name : zkx2024
// Author       : Jlan
// Email        : 15533610762@163.com
// Create Time  : 2024-07-31
// File Name    : const_tab.sv
// Module Name  :
// Called By    :
// Abstract     :
//
// 
// *********************************************************************************
// Modification History:
// Date         By              Version                 Change Description
// -----------------------------------------------------------------------
// 2024-07-31    Macro           1.0                     Original
//  
// *********************************************************************************
`ifndef  CONST_TAB 
`define  CONST_TAB

module const_tab #(
    parameter   W = 16
)(
    input   clk,
    input   rst_n,
    input   [8:0]   a,
    input   en,
    output logic    [2*W+1:0]   const_tab_out
);

logic   [47:0] cos_sin_out;

always_comb begin
   unique case(a[5:0])
        0:   const_tab_out = {24'd8387976, 24'd102941};
        1:   const_tab_out = {24'd8386081, 24'd205866};
        2:   const_tab_out = {24'd8382923, 24'd308761};
        3:   const_tab_out = {24'd8378503, 24'd411609};
        4:   const_tab_out = {24'd8372821, 24'd514395};
        5:   const_tab_out = {24'd8365878, 24'd617104};
        6:   const_tab_out = {24'd8357675, 24'd719720};
        7:   const_tab_out = {24'd8348214, 24'd822227};
        8:   const_tab_out = {24'd8337495, 24'd924610};
        9:   const_tab_out = {24'd8325521, 24'd1026855};
        10:   const_tab_out = {24'd8312293, 24'd1128944};
        11:   const_tab_out = {24'd8297813, 24'd1230864};
        12:   const_tab_out = {24'd8282084, 24'd1332598};
        13:   const_tab_out = {24'd8265107, 24'd1434132};
        14:   const_tab_out = {24'd8246886, 24'd1535449};
        15:   const_tab_out = {24'd8227423, 24'd1636536};
        16:   const_tab_out = {24'd8206720, 24'd1737376};
        17:   const_tab_out = {24'd8184782, 24'd1837954};
        18:   const_tab_out = {24'd8161611, 24'd1938255};
        19:   const_tab_out = {24'd8137211, 24'd2038265};
        20:   const_tab_out = {24'd8111586, 24'd2137968};
        21:   const_tab_out = {24'd8084739, 24'd2237348};
        22:   const_tab_out = {24'd8056675, 24'd2336392};
        23:   const_tab_out = {24'd8027397, 24'd2435084};
        24:   const_tab_out = {24'd7996910, 24'd2533409};
        25:   const_tab_out = {24'd7965219, 24'd2631353};
        26:   const_tab_out = {24'd7932329, 24'd2728900};
        27:   const_tab_out = {24'd7898244, 24'd2826036};
        28:   const_tab_out = {24'd7862969, 24'd2922747};
        29:   const_tab_out = {24'd7826510, 24'd3019018};
        30:   const_tab_out = {24'd7788873, 24'd3114834};
        31:   const_tab_out = {24'd7750063, 24'd3210181};
        32:   const_tab_out = {24'd7710085, 24'd3305044};
        33:   const_tab_out = {24'd7668947, 24'd3399410};
        34:   const_tab_out = {24'd7626653, 24'd3493264};
        35:   const_tab_out = {24'd7583211, 24'd3586592};
        36:   const_tab_out = {24'd7538627, 24'd3679379};
        37:   const_tab_out = {24'd7492908, 24'd3771613};
        38:   const_tab_out = {24'd7446060, 24'd3863278};
        39:   const_tab_out = {24'd7398091, 24'd3954362};
        40:   const_tab_out = {24'd7349008, 24'd4044850};
        41:   const_tab_out = {24'd7298818, 24'd4134729};
        42:   const_tab_out = {24'd7247529, 24'd4223986};
        43:   const_tab_out = {24'd7195149, 24'd4312606};
        44:   const_tab_out = {24'd7141684, 24'd4400577};
        45:   const_tab_out = {24'd7087145, 24'd4487885};
        46:   const_tab_out = {24'd7031538, 24'd4574517};
        47:   const_tab_out = {24'd6974872, 24'd4660460};
        48:   const_tab_out = {24'd6917156, 24'd4745702};
        49:   const_tab_out = {24'd6858398, 24'd4830229};
        50:   const_tab_out = {24'd6798607, 24'd4914028};
        51:   const_tab_out = {24'd6737793, 24'd4997087};
        52:   const_tab_out = {24'd6675963, 24'd5079394};
        53:   const_tab_out = {24'd6613129, 24'd5160936};
        54:   const_tab_out = {24'd6549298, 24'd5241701};
        55:   const_tab_out = {24'd6484481, 24'd5321676};
        56:   const_tab_out = {24'd6418688, 24'd5400850};
        57:   const_tab_out = {24'd6351928, 24'd5479210};
        58:   const_tab_out = {24'd6284211, 24'd5556746};
        59:   const_tab_out = {24'd6215548, 24'd5633444};
        60:   const_tab_out = {24'd6145949, 24'd5709294};
        61:   const_tab_out = {24'd6075424, 24'd5784285};
        62:   const_tab_out = {24'd6003985, 24'd5858404};
        63:   const_tab_out = {24'd5931641, 24'd5931641};
    endcase
end
logic   [47:0]  ham_win_512_out;

always_comb begin

   unique case(a[6:0])
        0: ham_win_512_out = { 24'd1342761, 24'd1342177};
        1: ham_win_512_out = { 24'd1347427, 24'd1344511};
        2: ham_win_512_out = { 24'd1356758, 24'd1351510};
        3: ham_win_512_out = { 24'd1370746, 24'd1363170};
        4: ham_win_512_out = { 24'd1389384, 24'd1379485};
        5: ham_win_512_out = { 24'd1412661, 24'd1400444};
        6: ham_win_512_out = { 24'd1440562, 24'd1426034};
        7: ham_win_512_out = { 24'd1473070, 24'd1456241};
        8: ham_win_512_out = { 24'd1510167, 24'd1491046};
        9: ham_win_512_out = { 24'd1551828, 24'd1530428};
        10: ham_win_512_out = { 24'd1598030, 24'd1574363};
        11: ham_win_512_out = { 24'd1648744, 24'd1622825};
        12: ham_win_512_out = { 24'd1703939, 24'd1675784};
        13: ham_win_512_out = { 24'd1763583, 24'd1733208};
        14: ham_win_512_out = { 24'd1827639, 24'd1795062};
        15: ham_win_512_out = { 24'd1896068, 24'd1861310};
        16: ham_win_512_out = { 24'd1968830, 24'd1931910};
        17: ham_win_512_out = { 24'd2045879, 24'd2006821};
        18: ham_win_512_out = { 24'd2127170, 24'd2085997};
        19: ham_win_512_out = { 24'd2212653, 24'd2169390};
        20: ham_win_512_out = { 24'd2302276, 24'd2256950};
        21: ham_win_512_out = { 24'd2395986, 24'd2348624};
        22: ham_win_512_out = { 24'd2493726, 24'd2444356};
        23: ham_win_512_out = { 24'd2595436, 24'd2544088};
        24: ham_win_512_out = { 24'd2701055, 24'd2647761};
        25: ham_win_512_out = { 24'd2810519, 24'd2755311};
        26: ham_win_512_out = { 24'd2923763, 24'd2866673};
        27: ham_win_512_out = { 24'd3040717, 24'd2981780};
        28: ham_win_512_out = { 24'd3161311, 24'd3100563};
        29: ham_win_512_out = { 24'd3285471, 24'd3222950};
        30: ham_win_512_out = { 24'd3413124, 24'd3348866};
        31: ham_win_512_out = { 24'd3544191, 24'd3478235};
        32: ham_win_512_out = { 24'd3678593, 24'd3610980};
        33: ham_win_512_out = { 24'd3816250, 24'd3747020};
        34: ham_win_512_out = { 24'd3957077, 24'd3886273};
        35: ham_win_512_out = { 24'd4100990, 24'd4028654};
        36: ham_win_512_out = { 24'd4247902, 24'd4174077};
        37: ham_win_512_out = { 24'd4397723, 24'd4322455};
        38: ham_win_512_out = { 24'd4550364, 24'd4473697};
        39: ham_win_512_out = { 24'd4705732, 24'd4627713};
        40: ham_win_512_out = { 24'd4863732, 24'd4784409};
        41: ham_win_512_out = { 24'd5024270, 24'd4943690};
        42: ham_win_512_out = { 24'd5187248, 24'd5105460};
        43: ham_win_512_out = { 24'd5352568, 24'd5269622};
        44: ham_win_512_out = { 24'd5520130, 24'd5436075};
        45: ham_win_512_out = { 24'd5689832, 24'd5604720};
        46: ham_win_512_out = { 24'd5861572, 24'd5775454};
        47: ham_win_512_out = { 24'd6035246, 24'd5948174};
        48: ham_win_512_out = { 24'd6210749, 24'd6122776};
        49: ham_win_512_out = { 24'd6387975, 24'd6299154};
        50: ham_win_512_out = { 24'd6566817, 24'd6477201};
        51: ham_win_512_out = { 24'd6747166, 24'd6656809};
        52: ham_win_512_out = { 24'd6928913, 24'd6837871};
        53: ham_win_512_out = { 24'd7111949, 24'd7020277};
        54: ham_win_512_out = { 24'd7296163, 24'd7203915};
        55: ham_win_512_out = { 24'd7481443, 24'd7388676};
        56: ham_win_512_out = { 24'd7667677, 24'd7574448};
        57: ham_win_512_out = { 24'd7854754, 24'd7761117};
        58: ham_win_512_out = { 24'd8042559, 24'd7948572};
        59: ham_win_512_out = { 24'd8230979, 24'd8136699};
        60: ham_win_512_out = { 24'd8419900, 24'd8325384};
        61: ham_win_512_out = { 24'd8609208, 24'd8514513};
        62: ham_win_512_out = { 24'd8798789, 24'd8703972};
        63: ham_win_512_out = { 24'd8988527, 24'd8893646};
        64: ham_win_512_out = { 24'd9178309, 24'd9083420};
        65: ham_win_512_out = { 24'd9368019, 24'd9273180};
        66: ham_win_512_out = { 24'd9557542, 24'd9462811};
        67: ham_win_512_out = { 24'd9746764, 24'd9652198};
        68: ham_win_512_out = { 24'd9935571, 24'd9841226};
        69: ham_win_512_out = { 24'd10123848, 24'd10029783};
        70: ham_win_512_out = { 24'd10311481, 24'd10217752};
        71: ham_win_512_out = { 24'd10498358, 24'd10405021};
        72: ham_win_512_out = { 24'd10684364, 24'd10591477};
        73: ham_win_512_out = { 24'd10869388, 24'd10777006};
        74: ham_win_512_out = { 24'd11053318, 24'd10961497};
        75: ham_win_512_out = { 24'd11236042, 24'd11144838};
        76: ham_win_512_out = { 24'd11417450, 24'd11326918};
        77: ham_win_512_out = { 24'd11597433, 24'd11507627};
        78: ham_win_512_out = { 24'd11775880, 24'd11686855};
        79: ham_win_512_out = { 24'd11952685, 24'd11864495};
        80: ham_win_512_out = { 24'd12127741, 24'd12040439};
        81: ham_win_512_out = { 24'd12300941, 24'd12214580};
        82: ham_win_512_out = { 24'd12472182, 24'd12386813};
        83: ham_win_512_out = { 24'd12641358, 24'd12557034};
        84: ham_win_512_out = { 24'd12808369, 24'd12725141};
        85: ham_win_512_out = { 24'd12973113, 24'd12891031};
        86: ham_win_512_out = { 24'd13135490, 24'd13054604};
        87: ham_win_512_out = { 24'd13295403, 24'd13215761};
        88: ham_win_512_out = { 24'd13452754, 24'd13374405};
        89: ham_win_512_out = { 24'd13607449, 24'd13530439};
        90: ham_win_512_out = { 24'd13759393, 24'd13683770};
        91: ham_win_512_out = { 24'd13908495, 24'd13834305};
        92: ham_win_512_out = { 24'd14054666, 24'd13981953};
        93: ham_win_512_out = { 24'd14197815, 24'd14126624};
        94: ham_win_512_out = { 24'd14337858, 24'd14268230};
        95: ham_win_512_out = { 24'd14474709, 24'd14406688};
        96: ham_win_512_out = { 24'd14608285, 24'd14541911};
        97: ham_win_512_out = { 24'd14738506, 24'd14673820};
        98: ham_win_512_out = { 24'd14865292, 24'd14802333};
        99: ham_win_512_out = { 24'd14988568, 24'd14927374};
        100: ham_win_512_out = { 24'd15108259 , 24'd15048866};
        101: ham_win_512_out = { 24'd15224292 , 24'd15166737};
        102: ham_win_512_out = { 24'd15336597 , 24'd15280915};
        103: ham_win_512_out = { 24'd15445106 , 24'd15391330};
        104: ham_win_512_out = { 24'd15549754 , 24'd15497917};
        105: ham_win_512_out = { 24'd15650477 , 24'd15600610};
        106: ham_win_512_out = { 24'd15747215 , 24'd15699348};
        107: ham_win_512_out = { 24'd15839908 , 24'd15794071};
        108: ham_win_512_out = { 24'd15928502 , 24'd15884721};
        109: ham_win_512_out = { 24'd16012941 , 24'd15971244};
        110: ham_win_512_out = { 24'd16093176 , 24'd16053587};
        111: ham_win_512_out = { 24'd16169158 , 24'd16131702};
        112: ham_win_512_out = { 24'd16240840 , 24'd16205539};
        113: ham_win_512_out = { 24'd16308180 , 24'd16275055};
        114: ham_win_512_out = { 24'd16371136 , 24'd16340208};
        115: ham_win_512_out = { 24'd16429671 , 24'd16400959};
        116: ham_win_512_out = { 24'd16483749 , 24'd16457269};
        117: ham_win_512_out = { 24'd16533338 , 24'd16509107};
        118: ham_win_512_out = { 24'd16578407 , 24'd16556439};
        119: ham_win_512_out = { 24'd16618930 , 24'd16599238};
        120: ham_win_512_out = { 24'd16654881 , 24'd16637478};
        121: ham_win_512_out = { 24'd16686239 , 24'd16671135};
        122: ham_win_512_out = { 24'd16712986 , 24'd16700190};
        123: ham_win_512_out = { 24'd16735104 , 24'd16724624};
        124: ham_win_512_out = { 24'd16752581 , 24'd16744423};
        125: ham_win_512_out = { 24'd16765405 , 24'd16759575};
        126: ham_win_512_out = { 24'd16773570 , 24'd16770070};
        127: ham_win_512_out = { 24'd16777070 , 24'd16775903};
        
   endcase
    
end 

wire [W-1:0] ham_win_512_out_ql = ham_win_512_out[23:0] >> (24-W);
wire [W-1:0] ham_win_512_out_qh = ham_win_512_out[47:24] >> (24-W);

always_ff @(posedge clk or negedge rst_n) begin
    if(!rst_n)begin
        const_tab_out   <= '0;
    end
    else if(en)
        casez(a[8:6])
            3'b000: const_tab_out   <= {1'b0,cos_sin_out[47:24],1'b0,cos_sin_out[23:0]};
            3'b01?: const_tab_out   <= {1'b0,ham_win_512_out_qh,1'b0,ham_win_512_out_ql};
            default: const_tab_out <= '0;
        endcase
end 
endmodule
`endif

